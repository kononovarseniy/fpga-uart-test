library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity UART is
	port (
		clk_i: in std_logic
		
		
	);
end entity;

architecture rtl of UART is
begin

end architecture;
